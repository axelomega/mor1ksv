`ifndef MOR1KX_SPRS_SVH
    `define MOR1KX_SPRS_SVH

    `define SPR_BASE(x)   (x/(2**11))
    `define SPR_OFFSET(x) (x%(2**11))

`endif
